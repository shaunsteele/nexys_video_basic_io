task basic_io_driver::do_drive();
    vif.drive(req.delay, req.buttons, req.switches);
endtask