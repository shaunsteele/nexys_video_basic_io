constraint c_cmd {cmd = UVM_WRITE || cmd = UVM_READ;}
