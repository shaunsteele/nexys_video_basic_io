// hvl_top.sv

module hvl_top;

import uvm_pkg::*;
import basic_io_test_lib_pkg::*;

initial begin
    run_test();
end

endmodule
