task axi_lite_driver::do_drive();
    vif.do_drive(req);
endtask
