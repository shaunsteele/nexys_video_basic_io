// top.sv

module top;

hvl_top();
hdl_top();

endmodule
