// basic_io_test_lib_pkg.sv

`include "uvm_macros.svh"

package basic_io_test_lib_pkg;

import uvm_pkg::*;

`include "basic_io_test_base.svh"
`include "basic_io_test.svh"

endpackage
