// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : tb
//
// File Name: axi_lite_monitor.sv
//
// Author   : Name   : Shaun Steele
//            Email  : shaun.steele.1020@gmail.com
//            Year   : 2025
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Wed Jan 29 00:00:49 2025
//=============================================================================
// Description: Monitor for axi_lite
//=============================================================================

`ifndef AXI_LITE_MONITOR_SV
`define AXI_LITE_MONITOR_SV

// You can insert code here by setting monitor_inc_before_class in file axi_lite.tpl

class axi_lite_monitor extends uvm_monitor;

  `uvm_component_utils(axi_lite_monitor)

  virtual axi_lite_bfm vif;

  axi_lite_config     m_config;

  uvm_analysis_port #(axi_lite_seq_item) analysis_port;

  axi_lite_seq_item m_trans;

  extern function new(string name, uvm_component parent);

  // Methods run_phase, and do_mon generated by setting monitor_inc in file axi_lite.tpl
  extern task run_phase(uvm_phase phase);
  extern task do_mon();

  // You can insert code here by setting monitor_inc_inside_class in file axi_lite.tpl

endclass : axi_lite_monitor 


function axi_lite_monitor::new(string name, uvm_component parent);
  super.new(name, parent);
  analysis_port = new("analysis_port", this);
endfunction : new


task axi_lite_monitor::run_phase(uvm_phase phase);
  `uvm_info(get_type_name(), "run_phase", UVM_HIGH)

  m_trans = axi_lite_seq_item::type_id::create("m_trans");
  do_mon();
endtask : run_phase


// Start of inlined include file tb/tb/include/axi_lite_do_mon.sv
task axi_lite_monitor::do_mon();
    forever @(posedge vif.clk)
    begin
        m_trans = axi_lite_seq_item::type_id::create("m_trans");
    end
endtask// End of inlined include file

// You can insert code here by setting monitor_inc_after_class in file axi_lite.tpl

`endif // AXI_LITE_MONITOR_SV

